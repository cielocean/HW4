//------------------------------------------------------------------------------
// Test harness validates hw4testbench by connecting it to various functional 
// or broken register files, and verifying that it correctly identifies each
//------------------------------------------------------------------------------

`include "regfile.v"

module hw4testbenchharness();

  wire[31:0]	ReadData1;	    // Data from first register read
  wire[31:0]	ReadData2;	    // Data from second register read
  wire[31:0]	WriteData;	    // Data to write to register
  wire[4:0]	  ReadRegister1;	// Address of first register to read
  wire[4:0]	  ReadRegister2;	// Address of second register to read
  wire[4:0]	  WriteRegister;  // Address of register to write
  wire		    RegWrite;	      // Enable writing of register when High
  wire		    Clk;		        // Clock (Positive Edge Triggered)

  reg         begintest;	// Set High to begin testing register file
  wire		    dutpassed;	// Indicates whether register file passed tests

  // Instantiate the register file being tested.  DUT = Device Under Test
  regfile DUT
  (
    .ReadData1(ReadData1),
    .ReadData2(ReadData2),
    .WriteData(WriteData),
    .ReadRegister1(ReadRegister1),
    .ReadRegister2(ReadRegister2),
    .WriteRegister(WriteRegister),
    .RegWrite(RegWrite),
    .Clk(Clk)
  );

  // Instantiate test bench to test the DUT
  hw4testbench tester
  (
    .begintest(begintest),
    .endtest(endtest), 
    .dutpassed(dutpassed),
    .ReadData1(ReadData1),
    .ReadData2(ReadData2),
    .WriteData(WriteData), 
    .ReadRegister1(ReadRegister1), 
    .ReadRegister2(ReadRegister2),
    .WriteRegister(WriteRegister),
    .RegWrite(RegWrite), 
    .Clk(Clk)
  );

  // Test harness asserts 'begintest' for 1000 time steps, starting at time 10
  initial begin
    begintest=0;
    #10;
    begintest=1;
    #1000;
  end

  // Display test results ('dutpassed' signal) once 'endtest' goes high
  always @(posedge endtest) begin
    $display("DUT passed?: %b", dutpassed);
  end

endmodule


//------------------------------------------------------------------------------
// Your HW4 test bench
//   Generates signals to drive register file and passes them back up one
//   layer to the test harness. This lets us plug in various working and
//   broken register files to test.
//
//   Once 'begintest' is asserted, begin testing the register file.
//   Once your test is conclusive, set 'dutpassed' appropriately and then
//   raise 'endtest'.
//------------------------------------------------------------------------------

module hw4testbench
(
// Test bench driver signal connections
input	   		  begintest,	// Triggers start of testing
output reg 		endtest,	// Raise once test completes
output reg 		dutpassed,	// Signal test result

// Register File DUT connections
input[31:0]		    ReadData1,
input[31:0]		    ReadData2,
output reg[31:0]	WriteData,
output reg[4:0]		ReadRegister1,
output reg[4:0]		ReadRegister2,
output reg[4:0]		WriteRegister,
output reg		    RegWrite,
output reg		    Clk
);

  // Initialize register driver signals
  initial begin
    WriteData=32'd0;
    ReadRegister1=5'd0;
    ReadRegister2=5'd0;
    WriteRegister=5'd0;
    RegWrite=0;
    Clk=0;
  end

  integer i;
  integer dec = 0;

  // Once 'begintest' is asserted, start running test cases
  always @(posedge begintest) begin
    endtest = 0;
    dutpassed = 1;
    #10


  // Test Case 1: 
  //   Write '42' to register 2, verify with Read Ports 1 and 2
  //   (Passes because example register file is hardwired to return 42)
  WriteRegister = 5'd2;
  WriteData = 32'd42;
  RegWrite = 1;
  ReadRegister1 = 5'd2;
  ReadRegister2 = 5'd2;
  #5 Clk=1; #5 Clk=0;	// Generate single clock pulse

  // Verify expectations and report test result
  if((ReadData1 != 42) || (ReadData2 != 42)) begin
    dutpassed = 0;	// Set to 'false' on failure
    $display("Test Case 1 Failed");
  end
  else begin
    $display("Test Case 1 Passed");
  end


  // Test Case 2: 
  //   Write '15' to register 2, verify with Read Ports 1 and 2
  //   (Fails with example register file, but should pass with yours)
  WriteRegister = 5'd2;
  WriteData = 32'd15;
  RegWrite = 1;
  ReadRegister1 = 5'd2;
  ReadRegister2 = 5'd2;
  #5 Clk=1; #5 Clk=0;

  if((ReadData1 != 15) || (ReadData2 != 15)) begin
    dutpassed = 0;
    $display("Test Case 2 Failed");
  end
  else begin
    $display("Test Case 2 Passed");
  end


  // Test Case 3:
  // Write Enable is broken / ignored – Register is always written to.
    WriteRegister = 5'd3;
    WriteData = 32'd20;
    RegWrite = 1; //should be disabled but broken
    ReadRegister1 = 5'd3;
    ReadRegister2 = 5'd3;
    #5 Clk=1; #5 Clk=0;

    if((ReadData1 != 20) || (ReadData2 != 20)) begin
      $display("Test Case 3 Passed (should fail)");
    end
    else begin
      dutpassed = 0;
      $display("Test Case 3 Failed (should fail): Write Enable is broken");
    end

  //Test Case 3.1: 
  // Test Write Enable (RegWrite)

  //write enable 1 to 0 (1 at test case 2)
  WriteRegister = 5'd2;
  WriteData = 32'd15;
  RegWrite = 0;
  ReadRegister1 = 5'd2;
  ReadRegister2 = 5'd2;
  #5 Clk=1; #5 Clk=0;

  if((ReadData1 != 15) || (ReadData2 != 15)) begin
    dutpassed = 0;
    $display("Test Case 3.1 Failed: regWrite (enable to disable) not working");
  end
  else begin
    $display("Test Case 3.1 Passed: regWrite (enable to disable) is working");
  end

  //write enable 0 to 1
  WriteRegister = 5'd2;
  WriteData = 32'd16;
  RegWrite = 0;
  ReadRegister1 = 5'd2;
  ReadRegister2 = 5'd2;
  #5 Clk=1; #5 Clk=0;

  if((ReadData1 != 16) || (ReadData2 != 16)) begin
    WriteRegister = 5'd2;
    WriteData = 32'd16;
    RegWrite = 1;
    ReadRegister1 = 5'd2;
    ReadRegister2 = 5'd2;
    #5 Clk=1; #5 Clk=0;

    if((ReadData1 != 16) || (ReadData2 != 16)) begin
      dutpassed = 0;
      $display("Test Case 3.1 Failed: regWrite (disable to enable) not working");
    end
    else begin
    $display("Test Case 3.1 Passed: regWrite (disable to enable) is working");
    end
  end
  
  // Test Case 4: 
  // Decoder is broken – All registers are written to

  //set all values to 25 (broken decoder)
  WriteData = 32'd25;
  RegWrite = 1;

  for (i=1; i<32; i = i+1) begin
    WriteRegister = i;
    #5 Clk=1; #5 Clk=0;
  end

  //reading values
  for (i=1; i<32; i = i+1) begin
    ReadRegister1 = i;
    ReadRegister2 = i;
    if((ReadData1 == 25) && (ReadData2 == 25)) begin
      dec = dec+1;
    end
  end

  if (dec == 31) begin
    $display("Test Case 4: registers 1-31 are set to 25");
  end

  // Test Case 4.1: 
  // Testing Decoder

  //set all register from 0-31 has been set to 25 (broken decoder)

//  generate
//    genvar i;
//     for (i=0; i<32; i = i+1) begin: writeregblk
//      WriteRegister = 5'di;
//      #5 Clk=1; #5 Clk=0;
//
//      if((ReadData1 != 15) || (ReadData2 != 15)) begin
//        dutpassed = 0;
//        $display("Test Case 4.1 Failed (setting all values to 15)");
//      end
//    end
//  endgenerate
  
  //set reg 31 to 16
  WriteRegister = 5'd31;
  WriteData = 32'd16;
  RegWrite = 1;
  ReadRegister1 = 5'd31;
  ReadRegister2 = 5'd31;
  #5 Clk=1; #5 Clk=0;

  RegWrite = 0; //disable regwrite
  //checking reg 31 value
  if((ReadData1 != 16) || (ReadData2 != 16)) begin
    dutpassed = 0;
    $display("Test Case 4.1 Failed: Decoder not working");
  end
  else begin
    //checking reg 1 to 30
    for (i=1; i<31; i = i+1) begin
      ReadRegister1 = i;
      ReadRegister2 = i;
      #5 Clk=1; #5 Clk=0;
      if((ReadData1 != 25) || (ReadData2 != 25)) begin
        dutpassed = 0;
        $display("Test Case 4.1 Failed: Decoder not working");
      end
    end
    $display("Test Case 4.1 Passed: Decoder is working");
  end


  // Test Case 5: 
  // Testing register 0
  // Should pass

  //setting register 0 to 15
  WriteRegister = 5'd0;
  WriteData = 32'd15;
  RegWrite = 1;
  ReadRegister1 = 5'd0;
  ReadRegister2 = 5'd0;
  #5 Clk=1; #5 Clk=0;

  //reads 0 
  if((ReadData1 != 0) || (ReadData2 != 0)) begin
    dutpassed = 0;
    $display("Test Case 5 Failed: register32zero not working");
  end
  //doesn't read 0 
  else begin
    $display("Test Case 5 Passed: register32zero is working");
  end


  // Test Case 6: 
  // Port 2 is broken and alawys reads register 17
  // Test case should fail
  WriteRegister = 5'd3;
  WriteData = 32'd10;
  RegWrite = 1;
  ReadRegister1 = 5'd3;
  ReadRegister2 = 5'd17;
  #5 Clk=1; #5 Clk=0;

  if(ReadData1 != ReadData2) begin
    dutpassed = 0;
    $display("Test Case 6 Failed (should fail): Port 1 and Port 2 read different registers");
  end
  else begin
    $display("Test Case 5 Passed (should fail): Port 1 and Port 2 read same register");
  end


  // All done!  Wait a moment and signal test completion.
  #5
  endtest = 1;

end

endmodule